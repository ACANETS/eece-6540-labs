��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-@���rahZ����*��:�>2/}nQ.��;�p� .��I��u�����c^�.���&��U�,<6V�/���i��?GQ�.��V��?oj�q��8}��	D���o ��Z�� �s�1c��K��ĘV�Z�~����p�l��?��R����lf-[W���f$�J�5��D:mb�@XNQT3�,�?F��3|�N4�����S �n/rq!�t�=�ohWt�_a�7|^���
��0���sW���IᡃEe!�`�(i38�I+�{�Ӓ���h����(Y��h_07��V��&|6�łZ��0y<j]��H]xGMG�2�3�0UhN%ׄ�ns6������y�2)��(p2p)'�8ϳ	}�e!��������߰��͠>��_���t��jo�eW-��ӓ'�al��paf��pD��<��3Z�a�²���C�V�^�"��J�"�퀢W�����*ú��ƞ�qx���J���֤X�j,Zs������gFUB;yB���x	�&"=G�H�D��Lh�&��?N�����Q���qa�EuK�}w�*�*���d����C1zh���
�]S:ֻ�K6ή-��8�#ohWt�_a�k�Ԧhg���'�al��p���B]5)�'�r��'q3�]qLC"{p�G��<��i�m���5�<��~A㉙��[6�)�}��K��;�/O�5'KL[���/*z+d�B�f��!�_��Ҿ��?�4�ʗ�m���;�L|�1��?�1˃�J\wu��v�<f)��,�c�|k�J��-�Y=�#��^ ���L�Y&ׇӭ��h��в���'͍�h\y ˊ�YN��{no�U��^*hrY���F1xH�#�rU҃��~��cC��O�-��8�� �k�IkY�G�
��L�矤�t:(�uO�v���S[W���;\=�H��CW\o6LԪ�u#7z�� Iô͚X?�o>�j��^ :��$q��mKx"E&��� ��l$�������-VLV,Z���ް��!����ˍ!`�^uf8�i�VK9�{F&�z��Iښ��}�2OŘ�C}���\�4�ʈK ������=�����Y�ۻp��@4�+h�	��ދ�*w��H�D�cBP���N�8�c�J���a\Y�����e��rט�������@Ő��t2(;����q�����d�0�YĊ���[ �����
���*,f$�7Q0- ��Ck�fÜ�2/���}������]�0�lK'���Xwʈ���m"p�ħƿ�9c�1��8�h����,����^�V�.��v'gn���1�/�Δ��IgPgud�����`UNP�V��o5]�t���Zu�Ì�s��X�e��ښ�s���I���b�⪒��S �=�[T�)�����5�VY(������b�Kzb�d&(C�#�7#^�Vn���4]�sV�"$�dg�ݚ�Н�:��9KmjWOPg��&yy�;�i*�f`�o�${U��w�X�|0����?�-� 
�FܔR'�Ϟ�Fa��ƙ�Q;��IjWOPg��&yy���͵���ݧG �ŴP��Cn�CIEn4];ˍH���]&�HF@��u�$�R�nl�;�w������4]�sV�"$�dg=wK��7�&7�ѐ�O2�;�
Q���n���i�H�yRN�]�5'�?�R+�{�!��_3#ڸZ鎬����op%�l�R�9����IN<��z��}�Q2�+�Y��
�q���:��{l�f|�ό���.Ӫm��k�p�|��].��'���Xw��4L2�����c-(��?()��Ä�'���Xw�!�Tc_j��r�.��:�W@�]�!����
u�P}W��_K����(�
t��Y�{'%s���'����-��qs�VYp��HM�e��`y����:M�'��,e(}���(�
t�ژq���U��>;8ψ`��L��s�|��].��'���Xw�j�7��o�${U��w�X�|0���ߪ��w��ѫ���;�.�xF���J�m��L�U�����>WԆ.l�~��X���]�!��UX���`���
�u:	�����Q0�b��&'�z��h��jg��ג&���?��A�����e�I����j���Q8� Lڈ�|��!n}y���q���U�9B36�CF?�(X��qp]3�އ�>���5iM�xq9g�M�G�n�Ѹ�(��c�27.l�G5�`�D3��E%�\��U@IE�U����S8�<�)��'��Q;��I��BT�^��a(􆿳�����|�z�ʵC<���}~q�K7G#+�Ǘ0z�cULh�K�}��h\���e�Q��'��j7�v�ԯ�`�L�i֭?�\���3cx���K*FX�H���@IE�U����S8���Z�/������i��BT�^��a(􆿳�����.q�<X��u�:l��Z+r��TD��ό���.�<��D�V�[�Gv��F��(�
t�ژq���U�(�v������6����Y�-�_{sx��(�
t�ژq���U��|ٚ�~�;�s�*�:�L��?�<O�����(�
t��Y�{'%s���'����-��qs�VYp��HM�e��`y������3'�L��1�G�Qc�k]m�����9�dMbZ鎬�������(����T�3,�t_-Z��T�\ �͆��X������XQ �Kk�2�"�z��"@IE�U��~j�9Y�=�����X����(h�š�b)��I�n�� Oag�qod�֓���X����(h�š�b)-�uA^�Ko�5����`K9g�M�G�n�؀���%Z鎬�������(���P�:ާ�zl���yp��HM�e�Nu�5=��l|�*"k��c��*��#�|.�Tӏ,b�-�lg�W8]��?|VO�⅘��]�!��	Ǹ�y85�b�S���}�0�7��65��
=k�� ��ł�!r�dN�<@Iv�����a�pzl��a��ӎ�Xp�,4�֧��L�q����f�:�ǯ��]�!��	Ǹ�y85��U�u��Za��Z���Ga(􆿳���Qs����I�O�D�P�_Q�����9�S��Y�Z鎬����Y�V��#q�������� f�Lu�m���H�p�'���Xwa'�<� \R?Jk`_>�Q�k^�ïw��O�$F�5�����'���Xwa'�<� \�㕀rW�*�u��6뎗0z�cULhv�R�+Z`�"�X��O�'{��T�\ ��}�of��zK��i�� La������t�f���L����]�!���1����m�9��׼���c-(��ܬ��x��!o�OB쓘q���U�pzl��a���-W?8B!��[u_ q1j�i��sD$���̷P��=�!��$Q�����/���4֋>a��\%�glg�W8]��?V�a�M����\��T��=��g��IC:��>(��怋j&6ְ1 ��ȉN*l)�}�����T��.��W����x�]�V��[�o��9���E�&����f��jv�!d*�[��T��ڏ�j�j]��n�hy�y4����V���I#���^�)�[#!��ᗾ��b� �k0�40�/�-�I�b�=fņ�a�t��Wgֲ lh�š�b)��)Ԙ+��ｗ��u��;e5V�]C��%��Ob���m��j#�{D�A�mJd���o��_�Rc0;�-��a���˗�
La���X!���*C���� ���{��W�����5d�B� ��~���4M̍���Qw�c4~Nrg�d�Z�X�#w��b܉�����	H5���ҡ}�%��v��jr�����c-(��ܬ��x��!I��Uo����\n0�8�&?ZX5����7`�5�o�������3��a���d�a@��n
V~$�M�Ki�Z�h��$�ð��TYeN�j�W�b܉�����	H5���ҡ}�]�[��*�mW[�Ƶ\����H�Ծ�6UQ�㔩�LA�dWH�:�g�"I��h;�ab���c-(��=��c���&?ZX5�I���H�گ���VPYUt�\�3H�f��OLa����R~k��d�ð��Tbݖq!��'�E�Jg�LA�dWH�:�g�"I'�^�����P�HS|�4�04�jf��Bǳ/i��f�iC���R~k��d�ð��T9��0'����f�iC������t�f����pD��=�<�^p�-a�D͢q��`�Lx(�i��/R#k�˟ܒ�o|k�Lb�5ߧE4��rw�&�z<a��N� φ��<�6��Q�zp���zj7i�j�9��Ң�M��;�	��}sc8��B���F�9g�M�G�n f�Lu�m��jЏ�_� f�Lu�mQ����`��'C�>��/����p��BZ��L(�0Q���g���C1zh9�n�p8hѶ���� f�Lu�m�� ���~�0Q���g
3K�������: a�`7�H'` �#����mW[�Ƶ\�ŋ~���%.ݒ�O�@C���� �u|Z�x��p����C�@^��}�/����p����E�i3���;���EWrC6�=�����!���w��z䮃������+U�HJ�hJ��Gݟ�����-VL�d�٣��c�A�L'��Av�Hѡ�\	��rR���"X��[N�f��*ތ+U�HJ�h2�}�Q�� ���˃�I�d�٣��c�A�L')6�Y������i�t_-Z��T�\ ��^*������;���EWrG9�:Q������M�q'���Xw�j�7��}M��+�.ީ �����owђN�~%鯅�����v�+�G���p� f�Lu�m�k]m���2$�q.e'���Xwd�n]N�P�:ާ�zl���yp��HM�e�Nu�5=��{=J���}�f��"�P�!�c��H>+�w�������+U�HJ�h�4zԞ7Y��0Y d���2$�q.e'���Xw{=J����$�,o��}�^<o}?Q2�+�Yɱg#����t|Ơ$��#8Ԧ�/#�c$?���rs�i���%��v���0�BE�9Y}��P���"X��[�`�L�i� ��b�FP&;w>`�2ݧ�&����<���՞e{*�u��6�Q2�+�Yɱg#������^�m����*6S�4��?��kR�KC�m��O*�u��6뎋�ġC��ׇ�������[�S�n�H[\�'��g�d��liJ�9J?#y�>�)L�*���ߡ|z�ä�@�Z��&61������m%�td7���{_8�Y��n3��v2���d2<��k]m��l|�*"k��͆�Wu"����S����(����D��Z�خ-�D��~4�ˇ�h��]�Hlu����C��!a/֐��̺�E�g������͆�Wu"�Z �I�Ӧ�}r�HDʞ�sB�_�����C���t:���Ϳ��RB�Wa/�o�@C��_��+������C�m�QA�Q* jr�����c-(����O� ��f;[���0���7�0>�Q�k^�ïw��O�$FP��{�/a�Mv!���xǦ"�7�F�Q�Y ����,��(p����c3����1j|g[Ҡ(Y�u�o���z!�l�����C�8$�*�J�Z���{lIk`��L��sE�g������c��*��#-���)��r��V�@�d��-��!���0I52znu4Bޗ����Lg�)I���H�������Ut�\��G=X���$�L݄䎒���F ���S�L�{Ut�\�P��S�~D���X'��o�$�0��d����1����_� f�Lu�mz���5|��j�;�����!q�����
�?<��{
��>��!DO&�k��Z�u f�Lu�m��1�_�5kM��}�H�$�|�K�g֓:lla�v�r��ɲ�ΥT�t��f�B��IȘ�i�E�����
�?<�v1a{J��`��Ks���x�ԉ�>�h�����#8Ԧ�/���= �#y�>�)L���:+Fwa�}?�N�*����4����Bf���rs�(�̴Y�{'%s��jb�ܳ�mT~1���n�����0Ezi�9��n ����TZ94�l9=�-"���pP�=��_��#*63�o��a0:���@ 2��ɛ�?ө0=�!�hj���*6S�4��?��kR�KC�m��Of�!���ٸ#P�j2E�?rn�U_����m��m������U%����f�=�(������5n�[�f���r���˃�I��$��g}g�W8]��?�Jw��3�c�}���Fo|k�Lb@Wh�q0���VW���a�D�$0�1����_� f�Lu�mz���5|��j�;�����!q�����
�?<��{
��>��!DO&�k��Z�u f�Lu�m��1�_�5�7<(�lb�<�䛄��\�e�E���Q'�z'٥��gV�L�2�r��Km�^6*�d7Ud��_Y1��X���yω��Hp9��Ǧ"�7�F�Q�Y ��+��8Щ�J����3QP�B�=sM�/>�9j]��n�hy����˦G�٥P5���rs�i��='̹Z�;PM �%�s���3D��T�c��o�${U��w�X�|0��r1U�%G��"L?���w35������/{�����Hp9���@�n~K�?�\���3cx���K*F��}v�R"�����C��$dM!3��� �r#�j�����'A^%�=�$.�h�6Q�7�Ԧ)�,�|^�����1g�W8]��?�̟�1��H�^W3����4��� {�'#��p�-a�D͢q��`�L�5ߧE4�� �U�O���iw�|�ݭ�̓u�J� f�Lu�m�k]m��?�qjv
Kð��T���cg�(����D��Z�خ-�D��~4�[8�[Kh���˃�IZ<��K�'���Xw�j�7����5�"�r����D��q&G��|n�W`�"�X��Nݲ���+��.�[ ٓ��r_��m�?�\���3cx���K*F��}v�R"m������ f�Lu�m�k]m��=�(����J�1����9�8;��Bǳ/i��f�iC���B�_�+�)1F#�֞q>l6� �	�ėX �����n]���� ��5�gZ���������>=�o*���=�7=���jV�w(��q4C��w��a�%L�`���žj)�����R�����G�h�`E�����-VL����v�?�����-VL'd��i�)<��D�V��*�V$ ��`��Ks���x�ԉ�>�%&^�nƒg�|R��q�q�����
�+���8�N]-?6���f�iC���B�_�+�)<���H;R�V|fėX ���G�U?�䍎a-6�Da�z�������omi7x��8fDd=ܙ`	��
-m/�k]m���Wa�>�q��k]m��}e�7�M�"�^���9f�vr2�����U��r�LH'�`0Q���g �^M0�yKm�G��5M�YYroEWuIDẋrB�R���>_��
-m/�k]m���Wa�>�q��k]m���D9De��w��a�%t�F]T 	��w��a�%��ЀFhxYeN�j�W��_��+������C�m�QA�Q* �K:+>. K ��XƤ5_�9g�M�G�nWKg�Vw_�Ut�\�0���7�0>�Q�k^��z�)A��j���x�ԉ�>T۳�͕��d�4�t��Է'�r��'q��{�������g�|R��qnX�i֝�x(�i��/R#k�˟ܒ�o|k�Lb_N���9��	���rFgK%qm�J+63�o��a0L>�v�{�WE� ��7ҩ���n
V~$���9���Q��v��u����)9�A��=ʻ������3gWaU �I�%�z�J��ސ�����nF���]�Hlu������:��KY�[b%Ɨ���|:w��!C���� ���ۀa��Ȭ�J���犩�I�9@'g���c%�%A��=ʻ������3�1ǺvK}��a-6�Da�Msc	�ۮ[�����a�vݝh�c�A�L'�n��ع��\���e�Q��e�p�^~>��m�"L?���M��ZLh-�� ���$�� ��6A��e-x�_�c�}���Fo|k�LbJ�1��슀.�[ ٓ��r_��m�ސ�����nF���]�Hlu���K���L����� +\�?��D�$0�	W��^$k���	HLS��Va�ir�a�Ho�ˆ�f#n�y�z�v嗏�iqI���
��D0^�!\����}r�HDʞ�sB�_��4y��ij-M�O��~�jr�����c-(����O� ����ΥT�t�L�.��ݾ9�d�L��Ӈ(j7h�A��	�_�z�T�D��r�:�
A*���ҍ緫ē!yX[�C����i������^`�|��K�z��KVY�/̥@X�4K%qm�J+63�o��a0��/S-�x{^4��*m e8�~��	W��^$k�6P�p�HZ#�+#��]#P�j2E�?T۳�͕��~��є27�C���� ���ۀa���u�1��s f�Lu�m�c5��c�}���Fo|k�Lb�"L?��ٶC$�-��k�����ش����-VL��(&y^,$X��WG ����L�ΪA�ʴ�!ޭđļw-b�&�I/��\]��a-6�Dajr�����c-(����O� ����ΥT�t�q�)]Q�x��r_��mjr�����c-(����O� ��+�AMm?��(xʶ���3*p�Hp�-a�D͢q��`�L�"L?��� e8�~��	W��^$k�6P�p�HZ~�똕<�/���jbPh79 ��/6�tTi���׏�����Mc�}���Fo|k�LbB�R���>_�/V�S���/���jbPhM�x���I�^A��x����
�?<I����P�J�1���K���L���4�04�jf&ظ����0o��,� f�Lu�mZU��<R �6��`��Q��v��u@�W`���joŶc0;�ļw-b�&�u�>Y�Ut�\���t6��ΥT�tB�R���>_lE��U���C��{/��K���L���4�04�jf&ظ���k�����ش����-VL��LG��&�h�6Q�7��ҿ�Gz��W ���tɣH���U����xQ�n
V~$0���7�0>�Q�k^�ïw��O�$FP��{�/a'٥��gV�T۳�͕��ɞJ$��^�5M�YYroE�4rh��|��3���ʪ���g�|R��qưb����+����,�x(�i��/RR���t�D�$0�`�|��K�zz��9�󔦵"�K�b��Ub�ۙD-M�O��~ӕ��d2<��k]m��������YC-�T^*��.�[ ٓ��4]a�#�b��nw;��-�?I�g��Q;��I�@�����Ut�\���"�oi�8+f«L�I�_Pg<˙Y�#�{U��"L?��ل��u
S�C�_]p���$�J�����u���^rYC-�T^*K���L���4�04�jf&ظ�����q\sv�I���и*�����x{^4��*m,�\����J���o3c�-��;���֤���n���v���=�W�� ����:+Fwa��˓#��͎>����'�r��'qm�±��m|/�l�`��\�806������X��֑xGV�z؝sK���L���4�04�jf&ظ���M���yt7�L8���q�n
V~$�Iw���L�8���-�r�MM�6�yJh�o�p�+���8ߏ[b%Ɨ�5%�h����v'#`�x��X��WG ���CnX�&��v~�z�xE�?F ����4D����'٥��gV�B�R���>_�S�V�C�d�����N���qHTZ_&bq�f;[���rw�&�z<a��r���#k�˟ܒ�o|k�Lb�%�`�ʾ@h����#o�]�ʄ�m�Թ���p�T��~��NC7�\��0׋e�4C�V�Q��3�� �f�˭�������VPYUt�\�����駈&����<���՞e{}�tJ�Ȫ��b܉�����	H5���ҡ}�6�+b�f� f�Lu�mz���5|� �O�)T۳�͕��`;��@�+;�6����O���H��`��Ks���ɛ�?ө�5ߧE4��rw�&�z<a.y�&5 �i�Y
�,�Ϭ��N��Y�#�{U�H\WC,߽��<�{~�1���'.5ko7�%���sC�CW�[��k�6o�d(�����lz�Q,~;�h�6Q�7� �^M0ܢ�$���45M�YYroEWuIDẋrG#��Ll(��?��kR�Ki�Y
�,˛AHCO�i�?��kR�KC�m��OK<桇d���_��+��
/<>��@"�^���9f�vr2�5ߥ�	K1�`�D3��暶/G��G9�:Q���i�֒�B�AKd��y c�󐪽�r���8��9�8,}'�%�y��A�����'�r��'q#�� �[N0�gŌa0�0Q���g
3K�������: a�`*l�\:6�
J���o3c�-��;��>�3�eZ~w����F�'�r��'qm�±��m|4��+$�P���(��[O��ɔ�<5���3��6?��[O��ɔ�<5���3��C�v��P�G=X��^M��C�\	��rR�c�3'A��0�7��65���KVY4n8�%�(%�ɏ�X,���֑xGV�05 S�s�l˛AHCO�i�?��kR�KC�m��O�|�vKSN���4]a�#�b��nw;��-�?I�g��Q;��I�@�����Ut�\�����
�?<���C1zhi�Y
�,x��F���kQ�Y ���|�vKSNҨ�(�l%�ɏ�X,���֑xGV�05 S�s�lrn�U_����m���yY�A1����
�?<�v1a{J�Ԧ)�,�|^�5ߧE4��}�)���x�ސ���ٰ�Ř�h�4M̍���it�V�Ԣ�Y9p��o��y��J*-M�O��~Ӊ�`�>`n-�b�F�F�Őue8�ސ�����H�^W3����4����Dr�2�}�u�0�_��/�ciJ�(?"��W����_�M86\�4�@����s��X��WG ����`�>`n-�b�F�F�Őue8�ސ�����H�^W3����4����Dr�2�p�-a�D͢fU�9�׏�����M��%�Lшφ��<�6�Ps_*�GqW�w��fD�B �n�6ӌ�Iۏ�.��]�xZPgud����;���O���)�l�n~��_eH�D���Lxx�rDcѴ��B�66��ѵ����j#�{D�A�mJd��K�����Ref/Лe�C�=���5�{4o-_j��r�.�h�!(C���� ��)h�j̎����F $u�ʹFJ�9o��;��
! R�7��1�G�Qc�k]m�����㺰�cC���� �]���5*_���g�|R��qưb�����_��hyM\�	8qLྫྷ��c\?
�����h	oS���\���l�©�}r�HDʞ�sB�_7s�9���of̲Az��%�g#����=��"��eer��,��]�!��	Ǹ�y85���~�S�8?��Z���Ga(􆿳���/�	1I��g#���rK��]�/p|VO�⅘��]�!��	Ǹ�y85�d�-�ð]�0�7��65��Wǖg3�MM
��,=^ħ(|`�Gu�#��nt�j�W���� ��;g�Y�{'%sgeߪ�{�e�X�+� �{�c�vI�ߪ��wQR�u9���+U�HJ�h<����y ����
�?<�v1a{J�ǃ4j�mrY�{'%s2�ew�n ����TZ94��owђN�~%鯅�����v�sk�TmU%����f�7s�9���of̲Az��%�g#�����!U�,�*�V$ �ǃ4j�mr�q���U�����v�y���jl7s�9���o@�ڗe' ��b�FP&x��F���kQ�Y ��*�u��6뎗0z�cUL�)��W�O��['����{:��$��a(􆿳��_����OO�;���EWr���1j|g[Ҡ(Y�u�o���z!�l7s�9���o@�ڗe' ��b�FP&���7��?�\���3cx���K*F��}v�R"7s�9���o 
���u N��r*a3�s�[a��vXٙZð��T��Ձm��J����FP?$�N(p����c3��z�������omi7x��8fDd=ܙ`	{�χI@�괆���-VL�ˇ�h��]�Hlu���E�Xf}}��v$���D�<D��-��r� DS�
�dN�<@Iv���a_|���x)��k\�7�ސ�����nF���]�Hlu����v�(�|�0Q���g �^M0�m�QA�Q* lE��U�����C�k�}��}N4����*��&�Hx��_�c�Z�~����v�� f�Lu�m̝' gi���Mv!���x�%&^�nƒg�|R��qưb�����|	ҷKD��ɛ�?өrn�U_����m��l|�*"k��͆�Wu"��@oX̥�2[O��ɔ�<5���3��< ���m�QA�Q* ��5n�[�f���r���˃�I��nF���-1QmO#��s��U;4@h����#o�]�ʄ�m�Թ���p�T��~���5|�d��G=X��{׳-�b���Ã�mH9��h��ۜ����KzMn
V~$���9���0Q���g	X��٤�Va�ir	�0��n�\�W�ECO�bԧLw�+�AMm?��D"x�A��,��5�Q	W��^$k�6P�p�HZN��6$��`ƺV���w35������C�ЋP����Hp9���@�n~K�?�\���3cx���K*F��}v�R"�����U��$dM!3��� �r#�j�����'����v�?MN*����$D\��z��@^��}�/����p����řA{��΄x�g��	��S8�'�}O[������Q����^kX��>ڑk��@ >t$���!���zl���y(ɹ�f=�>je`��@d:�����{~\�e�E���Q'�z�Mv!���xL�2�r��Km�^6*�d7Ud��_Y1��X�Jh�o�p��Hp9��Ǧ"�7�F�Q�Y ��b�� 4��P�!�c�dN��B���t^deZ���{lIk`��L��s�Y*&m1/��f���r8,}'�%�y�P�HS|�4�04�jfJߜ{�� ���aR��9�d�L�	�0��n�\�W�ECO�bԧLw�+�AMm?��D"x�A��,��5�Q	W��^$k�6P�p�HZy�&S��n�����؇0/���u
S�P�!�c�t}n�<�� #P�j2E�?fY�J�]�d(����D��Z�خ-�D��~4p��T�����$�����P�\�2����`jS������S�CП��/�����ྫྷ��c\?
������bR�Qa�vݝh�c�A�L'��Wm͏�rS�b�8Z�/����p���+=��B�n ����TZ94�l9=�-"���pP�=��_��#*63�o��a0:���@ 2��ɛ�?ө0=�!�hj���*6S�4��?��kR�KC�m��Of�!���ٸ#P�j2E�?rn�U_����m��m������U%����f�=�(������5n�[�f���r���˃�I��$��g}g�W8]��?�Jw��3�c�}���Fo|k�Lbx(�i��/R���3 ���|:w��!C���� ���ۀa��Ȭ�J����1���]]Q-�b�F�F����Y�/"�ސ�����@�`�\�e�E�~*�<�[�4b�-fz^)�hܮ��F�]؇��%��Ǐ�s|z�ä�@�Z��&61��T1�M�eer��,�������b'�Y@%��A<=ж<y�׀%\��������yω��Hp9��C6�=�����!���&v4�<0��.�[ ٓ�>1�8IpC���� ���ۀa��������tg?>l6� �	�ėX ��т1/�4o��Ut�\�������m%�td7���{_8�Y��n3��v2�@���J����p���$�J����3QP�B�=s�h�6Q�7��ҿ�Gz���D��B�UX���e��}r�HDʞ�sB�_�m����s�'�r��'qO�f
���"L?����@���J����p���$�J����3QP�B�=s�z�������omi7x�z����O'攤���}e�7�M�"�^���9f�vr2�����C�+/�����#�i�+?�|���˃�I)�>�$�>l�!q7��{n
V~$ɞJ$��^�5M�YYroEΖ�1�!�f'٥��gV�B�R���>_�����x�����Xf ��zR��%�>.}2�X>�Q�k^��vZ� �/Q(J�1���K���L���4�04�jf&ظ���U̿�n�5Km�^6*�d7Ud��_Y1��X�[Tj�qM�x3�ӬL��,�\�����\�W�EC�2[QvA��>�q��J|�����@CF���(٥P5���rs�i�̚irZ%���A+b���g�K�
�8���.�J��iU�ԝ5����pP�DI�-cv$���D�<D��-��r� DS�
���[Q���d7Ud��_Y1��X�O-�4'h��5ߧE4��@���i~ly	���rFgK%qm�J+63�o��a0L>�v�{�WE� ��7ҩ���n
V~$���9���Q��v��u����)9�A��=ʻ������3gWaU �I�%�z�J��ސ�����nF���]�Hlu������:��KY�[b%Ɨ���|:w��!C���� ���ۀa��Ȭ�J���犩�I�9@'g���c%�%A��=ʻ������3�1ǺvK}��a-6�Da�Msc	�ۮ[�����a�vݝh�c�A�L'�n��ع��\���e�Q��e�p�^~>��m�"L?���M��ZLh-�� ���$�� ��6A��e-x�_�c�}���Fo|k�LbJ�1��슀.�[ ٓ��r_��m�ސ�����nF���]�Hlu���K���L����� +\�?��D�$0�	W��^$k�&�c"�nU�[�ͬ�*�>WԆ.l&xPn�J1�̔��֤Z�h��ۜ��I�+�������:����XN˰Z�)&�}�Ȥ���n
V~$=�	�:˳����
�?<s��WM����x�ԉ�>���F��;Mݿ�N�\���I`��y�<zQ��������b9���<|���L�ΪA���XJ�;��zl���yM�0	�-1�g���ޔ7z�j�B�l<�䛄��=8{�u�>P�!�c��j$���X��WG ��~��є27�C���� ���ۀa���n��뾦��tTi����[b%Ɨ�jr�����c-(����O� ��+�AMm?��(xʶ���3*p�Hrw�&�z<a��r���T۳�͕��9�d�L�]c
j���ZVv ?Jѕh�蕡rUt�\��D�$0�\�e�E�0Hl&p?�ð��Th�Qf�=�	�:˳����
�?<s��WM����x�ԉ�>���pP�h�Qf�=�	�:˳����
�?<���z`��k��f�iC���B�_�+�)#P�j2E�?J�1���#P�j2E�?T۳�͕��~��є27�C���� ���ۀa���u�1��s f�Lu�m�c5��c�}���Fo|k�Lbrw�&�z<a��r�����˓#�������v�� f�Lu�m̝' gi��	W��^$k�6P�p�HZ�		�<�x�5ߧE4��p�-a�D͢q��`�L��/�ciJ��%�2X��<�(xʶ���,������P>l6� �	�ėX �����n]���\�e�E�0Hl&p?�U�.P	HȆ�:�M��f�Dj��UFe��x�ԉ�>��˓#���őT�ZS��A��H��p�-a�D͢q��`�L��/�ciJ�]c
j���\��buL���j���_��+������C�#o�]�ʄǚfA/kIIV�Q���a-6�DaC6�=�����!���P��
���A�)E��q�+���8ߏ[b%Ɨ��%&^�nƒg�|R��qưb�������VWO�}r�HDʞ�sB�_��F�İ���i����w:䩒=]'���3 ���}��0�g���ޔC�u�J�X\���e�Q^�;_�E�n
V~$��ӁW�^eer��,�NtZ��\���Jw��3��X�H��k��TA�l�Lɼ���t��3�*�I��f�^S�l�����z�/���
����~��&���j�W���?E�!$6�T۳�͕��{�χI@�괆���-VL����v�?�����-VLS��Õ��Jw��3�p�-a�D͢q��`�L��/�ciJ�"���u��A/�W�$�o�K�W��X��WG ��a�;�f����X��֑xGV�z؝s�l)�����k]m����.�[ ٓ��r_��m!s"֛
.C���~���J�������4�Ȭ�ӎ�Xp�,4�֧��L�q����*Y�Pܞ\p�-a�D͢q��`�L��/�ciJ�� ��5�gZ%�X�.���a-6�Da���1j|g[Ҡ(Y�u�o���z!�l�����C�&����1�6���f���˭�������VPYUt�\��Iw���L�8���-�r�MM�6�y��yω��Hp9����˓#���`;��@�+;�6����O���H��`��Ks���ɛ�?өx(�i��/R�-%��ʦ0rw�&�z<al����HZ� �U�O���5ߧE4��&��܏��O�͚��"�W�� ���*6�"�sC�CW�[��Q�
ֺ��⦚�%�4l�q#R���Z۳
0.P��{�/a�r-����g�y�ޥ-ju�u[�z�� �]	�c�C6�=�����!���5�<t]Y"�v$���D�<D��-��rv�V����v$���D�<D��-��r{R�@Mvu�>����9��0Y d���P�7ִ��#"�dN��B�y�J�#z�P�!�c��${`�J����#����p����B;�a��M��z����8�@ؾ�X��%&^�nƒg�|R��qu�V�D/����$���45M�YYroE�4rh��|�w�g�o�>����'�r��'qm�±��m|������E
! R�7��1�G�Qc�k]m���+��:H��
���׮w�v~�z�xE�?F �������p���v~�z�xE�?F ����=�(����|�'Ά��K3��N�r<���-,��n ����TZ94�7z�j�B�l�E8��5�:�Gé�ĻP�q����v�V����v$���D�<D��-��r{R�@Mv��a�z6�3��N�r<���-,��}M��+�.ީ ����7z�j�B�l�E8��5�:�Gé�ĻP�q����v�V���毾�P�\�2���?-Sah�"L?��٢p��vS���Dsw��J����� ʨ2X�P�!�cʍ����粧�?�\���3cx���K*F��}v�R"�ݾ-/̡#{W��:ԵưT҃�"�ޥG�@��UN����{^���2r0b�wa�����4��aa��x��Ut�\�?̝�7�䱟Bk���p?iAu�9���0��s��@^��}�/����p���x&n}(:W�6/�%��.T�����mz��c� �@w���H��j�Ï��	�M��.�X��a-6�Da?̝�7�䱟Bk���p?iAu�9���0��s��@^��}�/����p���x&n}(:Wx(�i��/RŻ�&ǥ���l0�Fi��|ր���5V��	��y9y�n&��J��<��%����<�k��m6[��e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc/?�s�m/C�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�yߪm����Y�{'%ssA'���?���ʢS����E@�ޗ9(����	�^��i�{���_�-h|,���(����>S��ә�����/�4�}n'���a*�x���� ��V�h����� ��?)��h�dZ�c��ǌM̯� VU+I���ť1k�`d��q�G����p��=.,����k����씧;�y������,�p���>��yܛ�	��|��	(���zL͊�q����N�:�Pn���������W;5B5Y+� �i7�sp>7.~Ƨ����?2^�9<o�nïi�JHn��z��r9�3/�OP�I^���V� D;5B5Y+�T�����N�܋�z2��~����ܷ|�p�6 �P�{n�da*;��;ۂ��IÙ=�H(c]9禩�5�Y�w��n	~����=��q�a\Y����_�G��GJHn��z���Z�n����t���i�Oa�b׉�^9Y�rU��6���h��J�1,!��a\Y����_�G��GJHn��z���YG�sT�Ș�TDв�0Z�׉�^9Y�rU��6���h�X��-�`V-u9�`�JHn��z���YG�s����Ӭ�oi�Oa�b�����I����ʮ�&3�-��_'��-d�Ry��\�v�[������ڶ�!!�+�R�G�Qr	�%\*��t���Y
 ����6?L���^ֻ����XP����d�ӓ
(~F�iO	������9`�p�0�B~W�u���iL�&Ш%� MjCЭ�J�1,!���i=���[&��?��
JHn��z���YG�s��K������-w˕��F��v_}*�����i��!�����9���k��h�@�sj|~��A�!`�u�!j;5B5Y+��q	k���Ak�$����v7�'��O�q�Yz��"�ձ[%�U��Q�f�!�+��7P��T�<��z��}�צ:�)��-��7�S�_�r-�Ճ)�E
Pv�~������]�!�����#ek�������:����7ѥ�"���$v�~������]�!�����#e;7mg�oc�.[K��m��/��*(�I�y.͸|��].��'���XwZ�֢t��FC5��v�c�.[K��m�u�M$S�{�,��TG���|���Aɘ%�ָkd�vu�Z��F����{l�f|�ό���.�2��T
�r��<Н?b���-(S�)37J*u.h�i�S�@����~��]��	B~��?b���-(S�)37J*u���
6��!l$P�ĝ�����-�$�<��z��}�Q2�+�Y��0]���!Vf����aU�7L�<��z��}拋ġC��ױ����h=�R��a:߻�%�q��{l�f|��rs�i���ZS��0���@	Q��"X��[?�e`N�aO'����M�{ET�\�%�OǱq�d�ֳ$7bOc� LҪ̏�7I�i����&���q�GR�c]�y����ҋX������S8�/��g��d\�p!|T����"X��[e�Xb��c���6�
y��i	3� ���ѡ�v�F#�5%� MjCИe��e�b]�lEGV`2B�7��MO���t�嗣H��BCk�2a�0/zﴚ�:�L��?�<O����!n}y��Y�{'%s�O��W��[�$��X�l�Lɼ�,0=]^	�&��������7LF��4�֧��L�q����[,��<5Z鎬�������(����|/��
3�b��nw;�X��������`y���e��~t�5M�YYroE�4rh��|��1�F�g�Z鎬�������l�T�|�1��?�WdM4@��2Smk0I��w��,c�A�L'�t�N)�~T-��qs�VY���/7R�%�T�\ ��U�f��4�tO��F'ot�k]m��8k>6s����]�!��	Ǹ�y85�ٙ�횔6�a\Y�����BT�^��a(􆿳�O�7�|lm�v|�ˑ����p|3�JR����TD���9�,�w�m����%�R/#٤M�i.�K�p}�����m/}|��XH�����,>$<�խ5�P�5�P3 C�0Q���g>y��d�,�Nn!���_��)�-pUO����LBTQ�C̱
^��%�a�������b�IeuѴ�8��ӳ�Y�
0������XP����|��{�r�\	��rR��y��O��톭��8h�U�$C�JrL�/H���H��߬���[>sd����MXݼ���jf&�~�7��MF�N�5pX�9��Ig`iZ鎬����D^Rm�	��f4!0v���=�%�1��w�&�=s9�E�m�b��곷Ї��u�\��~�A���Q�N�]�!���1����m�ρ;C���]����ڙc�К�^W�d�٣�����6>��b02�O �+s�ɔ�DY|5-��Y�Q3U�eT(�q���U�pzl��a��&5�/h�t���(�x��V����2B}G�J�ό���.�KX�U~�?E��T�ij�;{����Sx�lޞ�ό���.���K�Q���lp��V�j:e�KD��=Y��_Q2�+�Y�5�e`��9ꇤAfN�lR�����iͩ�;���Z鎬����Z��C�Ջ�n�\l����-~�*�[B�����'���Xw�j�7��ӣ��\g��@%:�����F1x
�ߴm�R�wX����K�Q��L�
�㱩� ���ﻋ-���C�M��N�۹t�������ͨk7����d��
F��=Y��_��ġC�����K�Qshf(�`�X�G[�Mf���9��Y�{'%s2�ew�}/A;T�c��iz�2��WX��y�g��U-�e5��e6²r,��>T�ї��;�
�{�4'��Xo��d޾ls'���Xwd�n]N�3g�Ƞ����i=���[�M*����9�ROe�Ё��������B�D�F ���>d��u�@}H�XC��k���4���>����Q2�+�Y�5�e`��9tteMh��v��'��e��"���N�_䈵vؐﻋ-���C�M��N�۔L�Xf1��V��&|6�łZ��0y#+�k�*�]�!���1����mr,��>T��pd����Y��'��e����9����@�f��l�q���U�pzl��a�x�-S����R��a�)�� ?ޏ'���Xwa'�<� \�]VI��Z/��������R��a�)�� ?ޏ'���Xwa'�<� \�&!�Tl�S� �D��>U�j����]�!���1����m���`�����f�����X�G[�M'�F2���ﻋ-���C�M��N��+w�7���[��:»}ю~VUo*��h9�'���Xwa'�<� \����9%=��M]l]�Qbi'D�ﻋ-���C�M��N���N��+�|�1��?�WdM4@Ȍ[PP�\��]�!��	Ǹ�y85�}�-���O��g���ޔ�h���o�8���/�a'�<� \�]VI��Za����g�cЉ�M��'ˑ�sO�rs�i�ק)"�僁Զ$�H� �b��nw;�X��������`y���pzl��a����������9�<��&�Rȧҟ�(((
�q���U�pzl��a��&5�/h�t���(�x�_S1�ޘ��]��K�ɿ�:8�cό���.���K�Q��p6Rh���>d���,f1P�y���O�.s�q���U�KX�U~�?���68�@�)��ї�!؈x.i����d�٣�����6>��r��&o�X�X�G[�

S{�M9�����O�w�&�T��>�%�*/��ġC���QK�>;?��Ϥk�;��|B}ø��y�w���H1��@�	��hN�q;�ǔ10\p c
N1�V&�����O�qTkή�Ádo�dvAg~�rk܀�#��˩���.|��f�ͣŗ�:���+"�9���B�I:׷�F�;�sB*�1v�!���y �谝��X�e�F����To?��m\Ӓ�qܛ�	��]���������ї4�z��pU6�M�S��2�{��΂IȀp/x��;�2V{D�G"�nT��z��uWU4y5=>F/�N��i+5�
�0�$�V�
�{�-靮a0r��:=�"ǭ{ �]�Kt�E*�#�,���ns)��E�$�v����ox3��vC��Z�G�a}Cy^6gV�+,:�� T<���^[ �1y�,	��"k@:G�	���=�ܾ�y�c��"x�O|?.����!��!����W�������9�xV��	7����G��O�L̍5��+'}����4L"�x��R�>(��F��eTQ�ȋ�V���w	����h _;��i�1�Q�^�� g�!�{5ܛ�	��A����¥��bMݪ��V�����׷eh��S�=�"�56RmHX���!���H���vO�[Jf퀔�������sr���0G3� B<���J��<��%����Y��EMܓ���;�e >���l�n�Zl�=%Fi]4�\��OA�z޷S�xo 7ǉ�&��8���������c-�z��~��D:<^��`Y�F�����I��<�|��F+��4���LT K���Db�J��@��$L��%��Z��b,7}��G���4��V*B�@,��ڬ�A ������ĎɌ�[9�-�Ҧ�{b�J��@��$L��%��Z��b,�0g���>a��v�<�RohWt�_a�fC��0��:Y����i%��ό�;�LȫԷ�/��Ϥk�;��|B}ø��y�w8#�RC�G�G~��6��YcN'�^������Q>�^2�����Vc2�����Vc2�����Vc�m7���e*bZ������&9����Ɵ�nKܦ��Fu)n2�����Vc2�����Vc2�����Vc͞����.�cF
'�q�f�_�oņ��>�䡓�1|��1y�HU����9/���`P�(r�7՚���[�V��j��R�`�7t}��ɬc��WNx�fr����_>V��@^0���'�$��S&ϊ��%�(j��yl�aY�`�8�N��2e�����'nZ/8G������ݨoa�I ����*�Z�s�ɞ�N6en-�@񔌞K�.%��s�)���_Zt�-MiЁ���0r�F�+�b�Ek�.��E����0��t:����I�n��!�P��l�s�f��ٸS|$vW�J^���[-���j��ku��s$y�t8ˎ8����A{�O�D)�A�� %�W�3ssc��w�,�Ǝ>c����2�AG�Ep��f&�Y;�t;z��r�B0�iY�<w&Rv 0��m#>�T�P��˳n1ja1�fT_UX��?bv�b��&J2�lt�E7���� X���������۞M�m:,�@���"~E��q8 r��!�W�,&��������}; ��`�V�F�P�_�^���\�}5�UI1�gB�� ]�Q%퇙?v���cc bާ�kU��*�E=w���������'|F������ґ�y�x$��ys\;��|B�˨Q{�(���t(&����2F����ӳ�Y�
�)�Ȍ�IP?�d���&�D�;E����.rV֡����=��|{� ��0h�5e�_c��p��S��ݬ"�b~*��s�F�KD�Vr[?z%CS2b�ү�+ҋj��)Ջ�z��"�����P��G�Q"���_ނMv!���x��%D�zQ��R��aI��%][��"��dr���L��Ń��$=��t���MIV��8Y��I/��\]��a-6�Da���[���8,b���-M�O��~Ӿ9�d�L���OW�+
դ>v��([��}qn
V~$�D�$0�x�-S����R��a�J��vT��N�g�c�` e8�~��m��"���@��b_їE���#P�j2E�?rn��<�ِmd���u�a��b<�C,�##P�j2E�?T۳�͕���{�Z՟|
[;T�!'ؔsy1�n��뾦� e8�~��5�UI1�gB�� ]�Q%�%��v�ڼtTi���׏�����M>je`��@d:�����{~��b����(K�Tl�;���f�����q9+t�}h�Qf�m��"���@��b�x�. ��#P�j2E�?�5ߧE4��c�}���Fo|k�Lbx(�i��/RŻ�&ǥ��a���F߸��S�Ȍ��"+VqS?�d���&��_WoI�Z4��=rf�\&�zI��������2F����ӳ�Y�
6:��d;��|Bp�%�Ut���w}�l�VH��T�<t��' ����X�G[�f׿�������!N�2��_:��y$[|�h���X ���ӳ�Y�
����.C؀(�2�x�X�!*�s����v`�9�PQ]�}K����M���(f���y���ri̲�=ީa)�!��ZB��,�Ӏ(�%�~3h���X �OLe�j�L�&�YڏR��!��ZB�ʳ87��Q�
#>:����0^��Q4K�Hk�t�迿��!�5m�)�T<��r)3nĉ�^P1~e�^jT����?e��g��A�i���g_mW�t���(�x��V���s_��!���j�s�PN�0O�4'��XoN���&��'��P��+BY��9�45��\1��jHM��Eؙ��?eY��5����G���:�?��V��h4���ӳ�Y�
����.C����>/�w-���V��&|6�łZ��0yI�[	ϱϲ�ΥT�tT۳�͕��rn��<�ِmd���u�a��b�g&xdp���ݾ-/���b練
��"�!�sp�	O�ƻ��W\D�F3���%Ff"�	-7���ү��d�<��7���n���&�Pݭ��%�x ~��O&�3�`�y�������"�X���G�����:�5Ӡ�X���e��
Ut�\�m��"���@��b�x�. ���s��U;4��:�E���[;T�!'ؔsy1�%��v��rw�&�z<a[5�M�����>d��u�@}H�XC��k���4Qa�D*O�amc�}�3�%Uo��� ��7CF��ܐ�}�S��/:+�e6j�"Hs�&_�f`��Zk��E�? +��^2�FP٫�]i�~,��.l��5'KL[��8�=w��imd��gޗ� �4A( 6�
�%{���܄��� M�=v��ۉ���o�TK������޷����"�<�6�Q=!X{�-i|�ZI��^���,f1P�y�VH��T�<�^~���QD9p;"��KO�#��K��%r]�Bа��Z�|>����wm�S� �D����a�Q��sH�}ˮ]ŧ��*
>2�dX�c���r�9��x�,f1P�y�VH��T�<�^~���QD���]���<�H�]����״P��l�GNj��	O�s�L�|[8�e�XC��yQ;�im���Lt���s��y$[|�h���X ��|��{�r�\	��rR�į������^�+�J�18].��@s��t:(ꚛ�[{i�����Ғ: ³s�Q;�m��~ж� ��%����p��B�Ա?�>����V;5h���X �����29��lӡ[L �$(r���3�k�� �9*���?�p~$J.r�J�}a>��V�!��ZB�*���d������OVe��˅�WR-���6Q��{�^�X�;٬sf.�T��T�ZT|�1��?�WdM4@�e��Y"��Q>�^2�����Vc2�����Vc2�����Vc ��xM��:@'�4��2~]��T?�7c��c��(ZH4~��2�����Vc2�����Vc2�����Vci�������]����ڙ�-�L�`�ح����7A�k�6��� ����ʕ�ӐDY|5-��Yb�58�D\�)�`"�:�>��g{n9�sn�X��̊�%�J)�h�O{�D~c*�y#�$?D�����:�3��~?ݤ�RD:9�ZM��#	�kW���������g��Z���CBZ�9����= �����D���5C�Z@e��3�!SC���H�8t�>�HcT�b�~G�e���巜j��fLe�]����>d���,f1P�ye��b���~�*�.i0/�]�s�����Rm)��%o��Pa�L��@X�h.P̐�R
�>������Yw��j�U�����GCc7�El����r0�N�������חo��� 3��H�̠��ç�B�;�y�>���/8'���/q�����v����oE.�q�2VP_ڍSSt�+F�'��,|RZ�YiD��Bd�Ҁv�i�K�%)3�d���P�f���>X�\m+Y�����!{��EFGbw�������a~bh?5膰�M�Ϩ<����p|3�z��a7��Q\9f��qb�Naْl��]�B}Ю�0U�L�#_���29a���Q������<�q}�w|�/U���!-�iP��G��\OL^��>%�Нo@���;1?�[F�sp֟kh�y��;��lMԲ���L��S-�����$þh���X �����R]Y�3�#�����T<�t�S�W���'h��� 5#�3֝��{�EG�'�fu��$lR�����i����)�j��dǑ؆�!��ZBU��<7�9�;��s\ڽS�����|�1��?���HEc-��0��"���
wh���X ���lp��f0{��
��8��E��Ia���F�笣�.Z;�������xa��rװ� t��]�qa]�݊3�m�E;���20ӠH��=w�A2ޮ}'�=��~6��_��jt0��Ƅ^�=�]�_Jz������D��ܒ0�=1E�Êp!!v*!��4�b�Eƃ��Q-s�b!��u���͂EC�y��Q28U�sQ��=d�Ɇ�X�$Z-�*�����-VL�z����9�j��f6&��?N����Sr� �A����ҹ��)U��XI��ׅy&�Zz�IÛ	���~��s��>�̔���c�(�3��[��\*n6�-�Ƙw���+t�a���`������w�=u�A��7X_��7��W`i�X�QK6�E����*��[�$��X�l�Lɼ���C�O�d�xǬa��u����9A���q�O�����¯�P��C	,��Ȃ�	�����'C`ø�X�t�G�����u�����&�܁�^����r
��Cݮ2�����sE���y1+�줥G��j�D�EH<J�B@��(�hS�}e�܍ˢO�bF_��a��Mz���O?�Sկw��[#M�4�!�["[:����!��lSԃ�0�!𨱹�I*�?��m�±��m|�Mpl�p�;�s�*�:�L�������-VL�++��Lm�>�Q�k^�ïw��O�$FOY�{�^��2��Z^��:���O�[a�vݝh�c�A�L'�8��Ns�[�$��X�/dΎ��^R�dm�Z鎬�������(����CTkd��a\Y���񺔗��FP�r�����L�
�T��i�e��F�2�\Ef�>���9x�=���&��^�,�<Zr���D�&x�Y���Q�@�<MN2��΢W&�]�רK̡g��b��y?����,\ަ�It*���1����nU��X|Qeu��<̐�<q�W��H/�/UMê�[�؀(�2�x@�����t��y�|�q���~�"����7Xa0~���;A���g�R�"i�g���h���R���ɢ���ڠ�Q;�m��j"^�����ϖ [@wPcIn-Hzn�!��ZB�;wJ��"tt�G�d�d�+��b2������ȼ�4�!O7I�"h#�)���w%e�D�m	$�WI��)A�
��v����=�\[L�R�X��Uq2��Z^��:�C�7�]���GljJ���a�X�� ��v|�ˑ����p|3�|6������:��;�jؾ�+Û�Dɰϐ�B��>����U:	��G���&���'b�'=�(W���\�����Vem.��;٬sf.��S�	�D��Og?6������p��U�)$���Ht��Չ�����l$P�ĝ��h�Q��p�ft��K<���q�� bާ�kU�������:�e9s�"�:7՟��"�]/���я�40��YS�k�� �9*���Q4uA����!Nǖ]��﹈�i�|54�
�ڧZ��7����.C����ꋖ��o��Ժ��e�����;��f��7ЋdU~���;AS�=hU�;�琾BT���h�}q~���Zy���4�e�e�{?�6�X�V��&|6�
#>:����0^���ז*��K*�lӡ[L ����h�}q���w�
Q0���ؽf���y3�/q�����;�
�{�4'��Xo�m,��"';�#��A	��e��Ż&3�-��_�Zl�<��?�d���&�D�;E��#�g��d�@���;�
�{�4'��Xo�,@� S�J �+s�ɔ��]����ڙ�k����ˇ�������r�G���Vem.�g��A�i�YW�S7�.����~j^�q�����f-(͕2�e(h0]�P��T��zw�\�ڧZ��7*M��J�<>�fpx���:�5Ӡ�q	�۝��&3�-��_��iz�2�nU>���g=��"�ԭd��g���V��&|6�łZ��0yI�[	ϱϲ�ΥT�tT۳�͕���w�����x0�Y��]&(K�Tl�;���f�����q9+t�}Ż�&ǥ��G^��w�&��E������;�
�{�4'��XoN���&��'��P��+BY��9�45��\1��jHM¸�k��CE]�٩��"�@�17ա1�\3�#j<��#����T���{�غŋ��6?L���x��y�o������w_	c��?:(?i˸3�J�
�M�'٥��gVا�˓#��͙�Og?6��m��"���@��b_їE����ݾ-/���b練��Og?6��z��"������@�a�ʢ�#vޖ�C�!��G�*s�D��	�LÉ7�tf�3�%Uo��� ��7CF��ܐ�}�S��/:+�e6j�"Hs<�?j=Ծ����dڐPSn��7i n�]|Y	@
�KS�'|�:w�`�w^���\�}+���Ã�&5�/hshf(�`�X�G[�{�[��/��5�P3 C��ґ�y�x��SrȎ�0h�5eו&��E������;�
�{�4'��XoN���&��'��P��+BY��9�:�d�~&3�-��_��iz�2�nU>���g=��"�ԭd��g���V��&|6�łZ��0yI�[	ϱϲ�ΥT�tT۳�͕���w�����x0�Y��]&(K�Tl�;���f�����q9+t�}Ż�&ǥ��G^��w�&��E������;�
�{�4'��XoN���&��'��P��+BY��9�:�d�~&3�-��_��iz�2�nU>���g=��"�ԭd��g��[;T�!'ؔsy1�n��뾦��"L?��٠����w_	c��?:(?i˸3�J�
�MɂMv!���x�5ߧE4��H��L�}wy�㱏>1�gB�� o� c ����D��n��2��F�0�ε�ތ�T>\��&�����bا*�W�Ǹ!2�͞nOY�c���ta���Om��g��%��&��p�h��в�������~�;|b[
.�sH�}ˮ�.���:\�� œ�Ę$����Z�g2*b���p6Rh���>d���,f1P�y�Ԡ�E���܄��� M��dW���݉�3�؞��&����,f1P�y�VH��T�<t��' ����X�G[Ἅ׉󾶓9�f?Y�O�Ķ�
�[�29a���Q�G���?�k�N�� �\	��rR�į������^�+�J��?��CG}	�Ճ��wqj��t���~���;AS�=hU�B����B��q.�)�l�do
<WAA �4A( 6'lg+������p߷Td��#��9@�;{�����%����	Q��|��RM����\(FK�T)O�K��:�g�@u^���ؽf��q.�)�l�dtO��F'ot�k]m���n��� �e����){���C�\Ef�>�77�qO!����C�/7���L>Q;�im���M:��2�n�ڤ���[U�&�n�����;���)�p*��PeD#���RDh���C�d��Iò҄;���[
�}3��*���1��²�=ީa)�!��ZB��,�Ӏ(��[��B�IxoҢbu�ߞ�(ɡ�>�(}%@��7�����fD�6:�Ӡ&F���x��az�d*�y3�/q��]Z3t<M`�ِ{o�7���B�=�7�V���үf�D=�
�a�� D��ﺣSq�#�-��>�C�~�)`� ��qQ��R��-���fx�Zq.�)�l�d �+s�ɔ�7�9���������D��h���_��Q�$G?q�a^z"�klʟ���Q��:'�T�r#�-m�f�����I A6˃rG%��/����&�h��(�5�P3 C��"r�V����U����BX�C����:�>��g{n9�sn�X��̊�%ę�Og?6�����lp�����2x^��x�e�w~U�I�cEY�����!{��E%���!j�_	c��?:(?i˸3���ޕa��W�\�9(xFog�[���V��ڧZ��7���%ݾ�8?�d���&�W����c�'��O�c%r]�Bа���/��D�jJ3�x0�Y��]&(K�Tl�;���f���� �z���@[�_zβrZ�tH�=��K�`�ν:qg�y��`';�#��A�V��&|6	��e��Ż&3�-��_�Zl�<��?�d���&�W����c�'��O�c%r]�Bа���/��D�jJ3�x0�Y��]&(K�Tl�;���f����Ps_*�GqW�w��fDk�F�ޗh�N��"���"�Y�%uрh�����;k�!!ʽ��?t�+)q�a^z"��v|�ˑ����p|3�|6������}[s��Wcu�5D��0h\Ef�>s�����g�0�u|x ����=f�����I A6˃rG�����<�4��:��v|�ˑ����p|3�l�1C��(��&5�/h�t���(�x�_S1�ޘ��]��Kоf�^P]W���g����/^�À<MN2��΢�9�2�L�t���(�x�_S1�ޘ��]��KЯ~ԫYc��LFC7�5$�)�vx�s��:��=VU�簦-�b�+�